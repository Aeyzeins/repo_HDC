module abc(

    input a,b,c
    output q
);


endmodule
