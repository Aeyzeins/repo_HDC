module example (
    input hi,
    output bye
);

    assign bye = hi;

endmodule
